`include "./adder.sv"

module cpu;

endmodule
